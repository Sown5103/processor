library verilog;
use verilog.vl_types.all;
entity signextend_vlg_vec_tst is
end signextend_vlg_vec_tst;
