library verilog;
use verilog.vl_types.all;
entity Mux21_32_vlg_vec_tst is
end Mux21_32_vlg_vec_tst;
