library verilog;
use verilog.vl_types.all;
entity AddSubtract_vlg_vec_tst is
end AddSubtract_vlg_vec_tst;
